class tx_sequence extends uvm_sequence #(tx_packet);
    `uvm_object_utils(tx_sequence)
    
    function new(string name = "tx_sequence");
        super.new(name);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        `uvm_info(get_type_name(), "Executing simple sequence", UVM_LOW)
    endfunction

    task pre_body();
        uvm_phase phase;
            `ifdef UVM_VERSION_1_2
            phase = get_starting_phase();
            `else
            phase = starting_phase;
            `endif
        if (phase != null) begin
            phase.raise_objection(this, get_type_name());
            `uvm_info(get_type_name(), "OBJECTION RAISED", UVM_MEDIUM)
        end
    endtask : pre_body

    task post_body();
        uvm_phase phase;
            `ifdef UVM_VERSION_1_2
            phase = get_starting_phase();
            `else
            phase = starting_phase;
            `endif
        if (phase != null) begin
            phase.drop_objection(this, get_type_name());
            `uvm_info(get_type_name(), "OBJECTION DROPPED", UVM_MEDIUM)
        end
    endtask : post_body
endclass


////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                         First Sequence                                   //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////



class simple_test extends tx_sequence;
    `uvm_object_utils(simple_test)

    function new (string name = "simple_test");
        super.new(name);
    endfunction

    task body();
        repeat(5) begin
            tx_packet pkt = tx_packet::type_id::create("pkt");
            start_item(pkt);
                pkt.randomize();
                `uvm_info("SEQ", $sformatf("Generate new item: %s", pkt.convert2str()), UVM_LOW)
      	    finish_item(pkt);
        end

    endtask
endclass   
class rx_sequence extends uvm_sequence#(rx_packet);
    `uvm_object_utils(rx_sequence)

    function new (string name = "rx_sequence");
    super.new(name);
    endfunction: new

    task pre_body();
        uvm_phase phase;
        `ifdef UVM_VERSION_1_2
            phase = get_starting_phase();
        `else
            phase = starting_phase;
        `endif
        if (phase != null) begin
            phase.raise_objection(this, get_type_name());
            `uvm_info(get_type_name(), "OBJECTION RAISED", UVM_MEDIUM)
        end
    endtask : pre_body

    task body();
        bit ok;
        set_response_queue_depth(-1);
    endtask: body

    task post_body();
        uvm_phase phase;
        `ifdef UVM_VERSION_1_2
            phase = get_starting_phase();
        `else
            phase = starting_phase;
        `endif
        if (phase != null) begin
            phase.drop_objection(this, get_type_name());
            `uvm_info(get_type_name(), "OBJECTION DROPPED", UVM_MEDIUM)
        end
    endtask : post_body

endclass: rx_sequence

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                          all_low                                          //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class all_low extends rx_sequence;
     `uvm_object_utils(all_low)

    function new (string name = "all_low");
        super.new(name);
    endfunction

    task body();
        //`uvm_info(get_type_name(), "Running all_low...", UVM_LOW)
        `uvm_do_with(req, {
            req.atready == 0;
            req.afvalid == 0;
            req.syncreq == 0;
            })
    endtask

endclass: all_low

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                      at_ready_high_only                                     //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class at_ready_high_only extends rx_sequence;
     `uvm_object_utils(at_ready_high_only)

    function new (string name = "at_ready_high_only");
        super.new(name);
    endfunction

    task body();
        //`uvm_info(get_type_name(), "Running at_ready_high_only...", UVM_LOW)
        `uvm_do_with(req, {
            req.atready == 1;
            req.afvalid == 0;
            req.syncreq == 0;
            })
    endtask

endclass: at_ready_high_only

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                          afvalid_high_only                                  //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class afvalid_high_only extends rx_sequence;
     `uvm_object_utils(afvalid_high_only)

    function new (string name = "afvalid_high_only");
        super.new(name);
    endfunction

    task body();
        //`uvm_info(get_type_name(), "Running afvalid_high_only...", UVM_LOW)
        `uvm_do_with(req, {
            req.atready == 0;
            req.afvalid == 1;
            req.syncreq == 0;
            })
    endtask

endclass: afvalid_high_only

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                          syncreq_high_only                                 //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class syncreq_high_only extends rx_sequence;
     `uvm_object_utils(afvalid_high_only)

    function new (string name = "syncreq_high_only");
        super.new(name);
    endfunction

    task body();
        `uvm_info(get_type_name(), "Running syncreq_high_only...", UVM_LOW)
        `uvm_do_with(req, {
            req.atready == 0;
            req.afvalid == 0;
            req.syncreq == 1;
            })
    endtask

endclass: syncreq_high_only

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                           rx_data_retention_seq                            //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class rx_data_retention_seq extends rx_sequence;
     `uvm_object_utils(rx_data_retention_seq)

    all_low low_seq;
    at_ready_high_only ready_seq;

    function new (string name = "rx_data_retention_seq");
        super.new(name);
    endfunction

    task body();
        `uvm_info(get_type_name(), "Running rx_data_retention_seq...", UVM_LOW)

        //Not receiving any atdata packet.
        repeat(20)
            `uvm_do(low_seq)
        
        
        //Here atready is 0
        repeat(5)
            `uvm_do(ready_seq)

    endtask

endclass: rx_data_retention_seq

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                           rx_flush_test_seq                                //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class rx_flush_test_seq extends rx_sequence;
     `uvm_object_utils(rx_flush_test_seq)

    all_low low_seq;
    at_ready_high_only ready_seq;
    afvalid_high_only valid_seq;

    function new (string name = "rx_flush_test_seq");
        super.new(name);
    endfunction

    task body();
        `uvm_info(get_type_name(), "Running rx_flush_test_seq...", UVM_LOW)

        //simple packet test, should recieve 15 full packets
        repeat(60)
            `uvm_do(ready_seq)

        //flush test, should receive 1 with atbytes = 3.
            `uvm_do(low_seq)
            `uvm_do(valid_seq)
            `uvm_do(ready_seq)

    endtask

endclass: rx_flush_test_seq


////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                           rx_ready_flag_seq                                //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class rx_ready_flag_seq extends rx_sequence;
     `uvm_object_utils(rx_ready_flag_seq)

    all_low low_seq;
    at_ready_high_only ready_seq;
    afvalid_high_only valid_seq;

    function new (string name = "rx_ready_flag_seq");
        super.new(name);
    endfunction

    task body();
        `uvm_info(get_type_name(), "Running rx_ready_flag_seq...", UVM_LOW)

        //Here atready is 1
        repeat(3)
            `uvm_do(ready_seq)
        
    endtask

endclass: rx_ready_flag_seq


////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                           rx_coherence_seq                                //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class rx_coherence_seq extends rx_sequence;
     `uvm_object_utils(rx_coherence_seq)

    at_ready_high_only ready_seq;
    
    function new (string name = "rx_coherence_seq");
        super.new(name);
    endfunction

    task body();
        `uvm_info(get_type_name(), "Running rx_coherence_seq...", UVM_LOW)

        repeat(32)
            `uvm_do(ready_seq)
        

    endtask

endclass: rx_coherence_seq


////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                           rx_byte_order_seq                                //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class rx_byte_order_seq extends rx_sequence;
     `uvm_object_utils(rx_byte_order_seq)

    at_ready_high_only ready_seq;
    
    function new (string name = "rx_byte_order_seq");
        super.new(name);
    endfunction

    task body();
        `uvm_info(get_type_name(), "Running rx_byte_order_seq...", UVM_LOW)

        repeat(40)
            `uvm_do(ready_seq)
        

    endtask

endclass: rx_byte_order_seq

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                           rx_valid_data_seq                                //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class rx_valid_data_seq extends rx_sequence;
     `uvm_object_utils(rx_valid_data_seq)

    all_low low_seq;
    at_ready_high_only ready_seq;
    afvalid_high_only valid_seq;
    
    function new (string name = "rx_valid_data_seq");
        super.new(name);
    endfunction

    task body();
        //`uvm_info(get_type_name(), "Running rx_valid_data_seq...", UVM_LOW)

        repeat(16) begin
            `uvm_do(ready_seq)
        end
        //     `uvm_do(valid_seq)
        //     //`uvm_do(valid_seq)
        //     `uvm_do(ready_seq)
        //    `uvm_do(low_seq)

    endtask

endclass: rx_valid_data_seq

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                           rx_at_bytes_seq                                //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class rx_at_bytes_seq extends rx_sequence;
     `uvm_object_utils(rx_at_bytes_seq)

    all_low low_seq;
    at_ready_high_only ready_seq;
    afvalid_high_only valid_seq;
    
    function new (string name = "rx_at_bytes_seq");
        super.new(name);
    endfunction

    task body();
        //`uvm_info(get_type_name(), "Running rx_at_bytes_seq...", UVM_LOW)

            repeat(25)
                `uvm_do(ready_seq)

            //atbytes 3
            // `uvm_do(low_seq)
            // `uvm_do(valid_seq)
            // `uvm_do(ready_seq)

            // `uvm_do(valid_seq)
            // `uvm_do(ready_seq)

            // `uvm_do(valid_seq)
            // `uvm_do(ready_seq)

    endtask

endclass: rx_at_bytes_seq

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////                         rx_exhaustive_seq                                  //////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

class rx_exhaustive_seq extends rx_sequence;
     `uvm_object_utils(rx_exhaustive_seq)

     at_ready_high_only ready_high;
     all_low            signals_low;
     afvalid_high_only  valid_seq;
    
    function new (string name = "rx_exhaustive_seq");
        super.new(name);
    endfunction

    task body();
        `uvm_info(get_type_name(), "Running rx_exhaustive_seq...", UVM_LOW)

         //simple packet test, should receive 250
        repeat(1000) 
            `uvm_do (ready_high)

        repeat(200)
            `uvm_do (signals_low)

        repeat(80)
         `uvm_do (ready_high)

        `uvm_do(signals_low)
        `uvm_do(valid_seq)
        `uvm_do(ready_high)
        
    endtask

endclass: rx_exhaustive_seq